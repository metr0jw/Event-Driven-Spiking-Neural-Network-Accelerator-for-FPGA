//-----------------------------------------------------------------------------
// Title         : Comprehensive Testbench for Synapse Array
// Project       : PYNQ-Z2 SNN Accelerator
// File          : tb_synapse_array.v
// Author        : Jiwoon Lee (@metr0jw)
// Description   : Rigorous verification of synapse array including:
//                 - Parallel BRAM banking
//                 - Weight configuration (single & batch)
//                 - Spike propagation accuracy
//                 - Timing verification
//                 - Stress testing
// Note          : Iverilog compatible version
//-----------------------------------------------------------------------------

`timescale 1ns / 1ps

module tb_synapse_array;

    //=========================================================================
    // Parameters
    //=========================================================================
    parameter NUM_AXONS         = 64;       // Scaled for simulation
    parameter NUM_NEURONS       = 64;
    parameter WEIGHT_WIDTH      = 8;
    parameter NUM_READ_PORTS    = 8;        // Parallel BRAM banks
    parameter AXON_ID_WIDTH     = $clog2(NUM_AXONS);
    parameter NEURON_ID_WIDTH   = $clog2(NUM_NEURONS);
    parameter USE_BRAM          = 1;
    parameter USE_DSP           = 1;
    
    parameter CLK_PERIOD        = 10;
    
    //=========================================================================
    // Signals
    //=========================================================================
    reg                         clk;
    reg                         rst_n;
    
    // Input spike interface
    reg                         spike_in_valid;
    reg [AXON_ID_WIDTH-1:0]     spike_in_axon_id;
    wire                        spike_in_ready;
    
    // Output spike interface
    wire                        spike_out_valid;
    wire [NEURON_ID_WIDTH-1:0]  spike_out_neuron_id;
    wire [WEIGHT_WIDTH-1:0]     spike_out_weight;
    wire                        spike_out_exc_inh;
    
    // Weight configuration interface
    reg                         weight_we;
    reg [AXON_ID_WIDTH-1:0]     weight_addr_axon;
    reg [NEURON_ID_WIDTH-1:0]   weight_addr_neuron;
    reg [WEIGHT_WIDTH:0]        weight_data;  // +1 for sign
    
    // Batch write interface
    reg                         batch_we;
    reg [AXON_ID_WIDTH-1:0]     batch_axon_id;
    reg [NUM_READ_PORTS*(WEIGHT_WIDTH+1)-1:0] batch_weights;
    reg [NEURON_ID_WIDTH-1:0]   batch_start_neuron;
    
    // Control & Status
    reg                         enable;
    wire                        busy;
    wire [31:0]                 spike_count;
    
    //=========================================================================
    // Test Statistics
    //=========================================================================
    integer test_num;
    integer test_passed;
    integer test_failed;
    integer output_count;
    integer total_output_count;
    integer i, j;
    
    // Expected outputs tracking
    reg [WEIGHT_WIDTH:0] expected_weight [0:NUM_NEURONS-1];
    reg [WEIGHT_WIDTH:0] received_weight [0:NUM_NEURONS-1];
    reg received_valid [0:NUM_NEURONS-1];
    
    //=========================================================================
    // DUT Instantiation
    //=========================================================================
    synapse_array #(
        .NUM_AXONS(NUM_AXONS),
        .NUM_NEURONS(NUM_NEURONS),
        .WEIGHT_WIDTH(WEIGHT_WIDTH),
        .NUM_READ_PORTS(NUM_READ_PORTS),
        .USE_BRAM(USE_BRAM),
        .USE_DSP(USE_DSP)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        
        .spike_in_valid(spike_in_valid),
        .spike_in_axon_id(spike_in_axon_id),
        .spike_in_ready(spike_in_ready),
        
        .spike_out_valid(spike_out_valid),
        .spike_out_neuron_id(spike_out_neuron_id),
        .spike_out_weight(spike_out_weight),
        .spike_out_exc_inh(spike_out_exc_inh),
        
        .weight_we(weight_we),
        .weight_addr_axon(weight_addr_axon),
        .weight_addr_neuron(weight_addr_neuron),
        .weight_data(weight_data),
        
        .batch_we(batch_we),
        .batch_axon_id(batch_axon_id),
        .batch_weights(batch_weights),
        .batch_start_neuron(batch_start_neuron),
        
        .enable(enable),
        .busy(busy),
        .spike_count(spike_count)
    );
    
    //=========================================================================
    // Clock Generation
    //=========================================================================
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end
    
    //=========================================================================
    // Output Monitor
    //=========================================================================
    always @(posedge clk) begin
        if (spike_out_valid) begin
            output_count <= output_count + 1;
            total_output_count <= total_output_count + 1;
            received_weight[spike_out_neuron_id] <= {spike_out_exc_inh, spike_out_weight};
            received_valid[spike_out_neuron_id] <= 1'b1;
            $display("  [%0t] Output: neuron=%0d, weight=%0d, exc_inh=%b",
                     $time, spike_out_neuron_id, spike_out_weight, spike_out_exc_inh);
        end
    end
    
    //=========================================================================
    // Tasks
    //=========================================================================
    task reset_dut;
        begin
            rst_n = 0;
            enable = 0;
            spike_in_valid = 0;
            spike_in_axon_id = 0;
            weight_we = 0;
            weight_addr_axon = 0;
            weight_addr_neuron = 0;
            weight_data = 0;
            batch_we = 0;
            batch_axon_id = 0;
            batch_weights = 0;
            batch_start_neuron = 0;
            output_count = 0;
            
            for (i = 0; i < NUM_NEURONS; i = i + 1) begin
                expected_weight[i] = 0;
                received_weight[i] = 0;
                received_valid[i] = 0;
            end
            
            #(CLK_PERIOD * 10);
            rst_n = 1;
            enable = 1;
            #(CLK_PERIOD * 5);
        end
    endtask
    
    task configure_weight_single;
        input [AXON_ID_WIDTH-1:0] axon_id;
        input [NEURON_ID_WIDTH-1:0] neuron_id;
        input [WEIGHT_WIDTH-1:0] weight;
        input exc_inh;
        begin
            @(posedge clk);
            weight_we <= 1;
            weight_addr_axon <= axon_id;
            weight_addr_neuron <= neuron_id;
            weight_data <= {exc_inh, weight};
            @(posedge clk);
            weight_we <= 0;
            #(CLK_PERIOD);
        end
    endtask
    
    task configure_weight_batch;
        input [AXON_ID_WIDTH-1:0] axon_id;
        input [NEURON_ID_WIDTH-1:0] start_neuron;
        input [NUM_READ_PORTS*(WEIGHT_WIDTH+1)-1:0] weights;
        begin
            @(posedge clk);
            batch_we <= 1;
            batch_axon_id <= axon_id;
            batch_start_neuron <= start_neuron;
            batch_weights <= weights;
            @(posedge clk);
            batch_we <= 0;
            #(CLK_PERIOD);
        end
    endtask
    
    task send_spike;
        input [AXON_ID_WIDTH-1:0] axon_id;
        begin
            @(posedge clk);
            spike_in_valid <= 1;
            spike_in_axon_id <= axon_id;
            
            // Wait for ready
            @(posedge clk);
            while (!spike_in_ready) @(posedge clk);
            
            spike_in_valid <= 0;
        end
    endtask
    
    task wait_idle;
        input integer extra_cycles;
        begin
            @(posedge clk);
            while (busy) @(posedge clk);
            repeat(extra_cycles) @(posedge clk);
        end
    endtask
    
    task clear_received;
        begin
            output_count = 0;
            for (i = 0; i < NUM_NEURONS; i = i + 1) begin
                received_weight[i] = 0;
                received_valid[i] = 0;
            end
        end
    endtask
    
    task run_test;
        input [256*8-1:0] test_name;
        begin
            test_num = test_num + 1;
            $display("\n=== Test %0d: %0s ===", test_num, test_name);
        end
    endtask
    
    task check_pass;
        input [256*8-1:0] msg;
        begin
            $display("  PASS: %0s", msg);
            test_passed = test_passed + 1;
        end
    endtask
    
    task check_fail;
        input [256*8-1:0] msg;
        begin
            $display("  FAIL: %0s", msg);
            test_failed = test_failed + 1;
        end
    endtask
    
    //=========================================================================
    // Test Cases
    //=========================================================================
    initial begin
        $display("===============================================");
        $display("  Synapse Array Comprehensive Testbench");
        $display("===============================================");
        $display("  NUM_AXONS: %0d", NUM_AXONS);
        $display("  NUM_NEURONS: %0d", NUM_NEURONS);
        $display("  NUM_READ_PORTS (BRAM Banks): %0d", NUM_READ_PORTS);
        $display("  USE_BRAM: %0d, USE_DSP: %0d", USE_BRAM, USE_DSP);
        $display("===============================================");
        
        test_num = 0;
        test_passed = 0;
        test_failed = 0;
        total_output_count = 0;
        
        //=====================================================================
        // Test 1: Basic Reset
        //=====================================================================
        run_test("Basic Reset Verification");
        reset_dut();
        if (spike_count == 0) check_pass("Spike count is zero after reset");
        else check_fail("Spike count not zero");
        
        if (!busy) check_pass("Array not busy after reset");
        else check_fail("Array busy after reset");
        
        if (spike_in_ready) check_pass("Ready to accept spikes");
        else check_fail("Not ready after reset");
        
        //=====================================================================
        // Test 2: Single Weight Configuration
        //=====================================================================
        run_test("Single Weight Configuration");
        reset_dut();
        
        // Configure weight for axon 0, neuron 0
        configure_weight_single(0, 0, 8'd100, 1'b1);
        configure_weight_single(0, 1, 8'd50, 1'b0);  // Inhibitory
        #(CLK_PERIOD * 10);
        
        check_pass("Weight configuration completed");
        
        //=====================================================================
        // Test 3: Single Spike Propagation
        //=====================================================================
        run_test("Single Spike Propagation");
        reset_dut();
        clear_received();
        
        // Configure some weights for axon 0
        for (i = 0; i < 8; i = i + 1) begin
            configure_weight_single(0, i[NEURON_ID_WIDTH-1:0], 8'd10 + i[7:0]*10, 1'b1);
        end
        
        #(CLK_PERIOD * 20);
        
        // Send spike from axon 0
        send_spike(0);
        wait_idle(200);
        
        $display("  Output count: %0d (expected >=8)", output_count);
        if (output_count >= 8) check_pass("Got expected outputs");
        else check_fail("Insufficient outputs");
        
        //=====================================================================
        // Test 4: Parallel Read Verification
        //=====================================================================
        run_test("Parallel Read (BRAM Banking)");
        reset_dut();
        clear_received();
        
        // Configure weights for all neurons from axon 1
        for (i = 0; i < NUM_NEURONS; i = i + 1) begin
            configure_weight_single(1, i[NEURON_ID_WIDTH-1:0], i[7:0], 1'b1);
        end
        
        #(CLK_PERIOD * 100);
        
        // Send spike and verify parallel output
        send_spike(1);
        wait_idle(300);
        
        $display("  All neurons received: %0d (expected %0d)", output_count, NUM_NEURONS);
        if (output_count == NUM_NEURONS) check_pass("All neurons received");
        else check_fail("Not all neurons received");
        
        //=====================================================================
        // Test 5: Inhibitory Weights
        //=====================================================================
        run_test("Inhibitory Weight Propagation");
        reset_dut();
        clear_received();
        
        // Configure mix of excitatory and inhibitory
        for (i = 0; i < NUM_NEURONS; i = i + 1) begin
            configure_weight_single(2, i[NEURON_ID_WIDTH-1:0], 8'd100, (i % 2) ? 1'b1 : 1'b0);
        end
        
        #(CLK_PERIOD * 100);
        
        send_spike(2);
        wait_idle(300);
        
        // Verify some inhibitory weights received
        if (output_count > 0) check_pass("Inhibitory weights propagated");
        else check_fail("No outputs");
        
        //=====================================================================
        // Test 6: Multiple Axon Spikes
        //=====================================================================
        run_test("Multiple Axon Sequential Spikes");
        reset_dut();
        clear_received();
        
        // Configure weights for multiple axons
        for (j = 0; j < 4; j = j + 1) begin
            for (i = 0; i < 8; i = i + 1) begin
                configure_weight_single(j[AXON_ID_WIDTH-1:0], i[NEURON_ID_WIDTH-1:0], (j * 16 + i), 1'b1);
            end
        end
        
        #(CLK_PERIOD * 100);
        
        // Send spikes from multiple axons
        send_spike(0);
        wait_idle(100);
        clear_received();
        
        send_spike(1);
        wait_idle(100);
        
        if (output_count > 0) check_pass("Multiple axons processed correctly");
        else check_fail("No output from second axon");
        
        //=====================================================================
        // Test 7: Busy Signal Verification
        //=====================================================================
        run_test("Busy Signal Verification");
        reset_dut();
        
        // Configure weights
        for (i = 0; i < NUM_NEURONS; i = i + 1) begin
            configure_weight_single(4, i[NEURON_ID_WIDTH-1:0], 8'd50, 1'b1);
        end
        
        #(CLK_PERIOD * 100);
        
        send_spike(4);
        
        // Check busy goes high
        #(CLK_PERIOD * 2);
        if (busy) check_pass("Busy signal asserted during processing");
        else check_fail("Busy signal not asserted");
        
        wait_idle(300);
        if (!busy) check_pass("Busy signal deasserted after completion");
        else check_fail("Busy signal stuck high");
        
        //=====================================================================
        // Test 8: Zero Weight Handling
        //=====================================================================
        run_test("Zero Weight Handling");
        reset_dut();
        clear_received();
        
        // Configure zero weights - should not produce output
        for (i = 0; i < NUM_NEURONS; i = i + 1) begin
            configure_weight_single(5, i[NEURON_ID_WIDTH-1:0], 8'd0, 1'b1);
        end
        
        #(CLK_PERIOD * 100);
        
        send_spike(5);
        wait_idle(300);
        
        // Zero weights should NOT produce outputs (filtered)
        $display("  Zero weight outputs: %0d", output_count);
        if (output_count == 0) check_pass("Zero weights filtered correctly");
        else check_fail("Zero weights should be filtered");
        
        //=====================================================================
        // Test 9: Maximum Weight
        //=====================================================================
        run_test("Maximum Weight Value");
        reset_dut();
        clear_received();
        
        configure_weight_single(6, 0, 8'hFF, 1'b1);  // Max weight
        
        #(CLK_PERIOD * 20);
        
        send_spike(6);
        wait_idle(200);
        
        if (received_weight[0] == {1'b1, 8'hFF}) check_pass("Max weight preserved");
        else begin
            $display("  Got: %h, Expected: %h", received_weight[0], {1'b1, 8'hFF});
            check_fail("Max weight not preserved");
        end
        
        //=====================================================================
        // Test 10: Last Axon Access
        //=====================================================================
        run_test("Last Axon ID Access");
        reset_dut();
        clear_received();
        
        // Configure weight for last axon
        configure_weight_single(NUM_AXONS-1, 0, 8'd123, 1'b1);
        
        #(CLK_PERIOD * 20);
        
        send_spike(NUM_AXONS-1);
        wait_idle(200);
        
        $display("  Last axon ID: %0d, outputs: %0d", NUM_AXONS-1, output_count);
        if (output_count > 0) check_pass("Last axon ID works");
        else check_fail("Last axon ID failed");
        
        //=====================================================================
        // Test 11: Last Neuron Access
        //=====================================================================
        run_test("Last Neuron ID Access");
        reset_dut();
        clear_received();
        
        configure_weight_single(7, NUM_NEURONS-1, 8'd77, 1'b1);
        
        #(CLK_PERIOD * 20);
        
        send_spike(7);
        wait_idle(200);
        
        $display("  Last neuron ID: %0d, valid: %0d", NUM_NEURONS-1, received_valid[NUM_NEURONS-1]);
        if (received_valid[NUM_NEURONS-1]) check_pass("Last neuron ID received");
        else check_fail("Last neuron ID not received");
        
        //=====================================================================
        // Test 12: Enable/Disable Control
        //=====================================================================
        run_test("Enable/Disable Control");
        reset_dut();
        clear_received();
        
        configure_weight_single(8, 0, 8'd100, 1'b1);
        #(CLK_PERIOD * 20);
        
        // Disable
        enable = 0;
        spike_in_valid = 1;
        spike_in_axon_id = 8;
        #(CLK_PERIOD * 50);
        spike_in_valid = 0;
        
        if (output_count == 0) check_pass("Disabled array produces no output");
        else check_fail("Output despite disabled");
        
        // Re-enable
        enable = 1;
        #(CLK_PERIOD * 10);
        
        //=====================================================================
        // Test 13: Spike Count Register
        //=====================================================================
        run_test("Spike Count Register");
        reset_dut();
        
        configure_weight_single(10, 0, 8'd50, 1'b1);
        #(CLK_PERIOD * 20);
        
        send_spike(10);
        wait_idle(100);
        send_spike(10);
        wait_idle(100);
        send_spike(10);
        wait_idle(100);
        
        $display("  Spike counter: %0d", spike_count);
        if (spike_count >= 3) check_pass("Spike counter accurate");
        else check_fail("Spike counter inaccurate");
        
        //=====================================================================
        // Summary
        //=====================================================================
        $display("\n===============================================");
        $display("  Test Summary");
        $display("===============================================");
        $display("  Total Tests: %0d", test_passed + test_failed);
        $display("  Passed: %0d", test_passed);
        $display("  Failed: %0d", test_failed);
        $display("  Total spikes processed: %0d", spike_count);
        $display("  Total outputs generated: %0d", total_output_count);
        $display("===============================================");
        
        if (test_failed == 0)
            $display("  ALL TESTS PASSED!");
        else
            $display("  SOME TESTS FAILED!");
        
        $display("===============================================\n");
        
        #(CLK_PERIOD * 10);
        $finish;
    end
    
    //=========================================================================
    // Waveform Dump
    //=========================================================================
    initial begin
        $dumpfile("tb_synapse_array.vcd");
        $dumpvars(0, tb_synapse_array);
    end
    
    //=========================================================================
    // Timeout
    //=========================================================================
    initial begin
        #(CLK_PERIOD * 500000);
        $display("ERROR: Simulation timeout!");
        $finish;
    end

endmodule
